module top_module( input a,b,c,output k,l,m,n );
    
    assign k = a; 
    assign l = b;
    assign m = b;
    assign n = c;
endmodule
